module c17(N1, N2, N3, N6, N7, N22, N23);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire _05_;
  input N1;
  wire N1;
  wire N10;
  wire N11;
  wire N16;
  wire N19;
  input N2;
  wire N2;
  output N22;
  wire N22;
  output N23;
  wire N23;
  input N3;
  wire N3;
  input N6;
  wire N6;
  input N7;
  wire N7;
  assign _00_ = N1 & N3;
  assign _01_ = N3 & N6;
  assign _02_ = N2 & N11;
  assign _03_ = N11 & N7;
  assign _04_ = N10 & N16;
  assign _05_ = N16 & N19;
  assign N22 = ~ _04_;
  assign N23 = ~ _05_;
  assign N10 = ~ _00_;
  assign N11 = ~ _01_;
  assign N16 = ~ _02_;
  assign N19 = ~ _03_;
endmodule