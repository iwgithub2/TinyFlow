module Mult(a, b, c
);
    assign c = a | b;

endmodule
