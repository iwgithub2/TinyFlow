{
  "library": {
    "name": "TinyLEF",
    "version": "1.0",
    "description": "Minimal LEF-style library"
  },
  "cells": {
    "NAND2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [8, 16, 10, 18] }
          ]
        },
      },
    },
    "MUX2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "s": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [8, 16, 10, 18] }
          ]
        },
      },
    },
    "AOI21D1": {
      "class": "CORE",
      "size": [30, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "b": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "z": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [8, 16, 10, 18] }
          ]
        },
      },
    },
    "XOR2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [8, 16, 10, 18] }
          ]
        },
      },
    },
    "INVD1": {
      "class": "CORE",
      "size": [10, 10],
      "pins": {
        "a": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "out": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [8, 16, 10, 18] }
          ]
        },
      },
    },
    "NOR2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [2, 6, 4, 8] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [8, 16, 10, 18] }
          ]
        },
      },
    }
  }
}