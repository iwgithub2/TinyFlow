
module TESTER (
  input clk,
  output reg unsigned data = 0
);

endmodule
