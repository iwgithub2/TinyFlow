{
  "library": {
    "name": "TinyLEF",
    "version": "1.0",
    "description": "Minimal LEF-style library"
  },
  "cells": {
    "NAND2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 7, 3, 9] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 3, 3, 5] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [12, 4, 14, 6] }
          ]
        }
      }
    },
    "MUX2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 7, 3, 9] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 3, 3, 5] }
          ]
        },
        "s": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 5, 3, 7] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [12, 4, 14, 6] }
          ]
        }
      }
    },
    "AOI21D1": {
      "class": "CORE",
      "size": [30, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 7, 3, 9] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 3, 3, 5] }
          ]
        },
        "b": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 5, 3, 7] }
          ]
        },
        "z": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [27, 4, 29, 6] }
          ]
        }
      }
    },
    "XOR2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 7, 3, 9] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 3, 3, 5] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [12, 4, 14, 6] }
          ]
        }
      }
    },
    "INVD1": {
      "class": "CORE",
      "size": [10, 10],
      "pins": {
        "a": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 4, 3, 6] }
          ]
        },
        "out": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [7, 4, 9, 6] }
          ]
        }
      }
    },
    "NOR2D1": {
      "class": "CORE",
      "size": [15, 10],
      "pins": {
        "a1": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 7, 3, 9] }
          ]
        },
        "a2": {
          "direction": "INPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [1, 3, 3, 5] }
          ]
        },
        "y": {
          "direction": "OUTPUT",
          "use": "SIGNAL",
          "ports": [
            { "layer": "M1", "rect": [12, 4, 14, 6] }
          ]
        }
      } 
    }
  }
}